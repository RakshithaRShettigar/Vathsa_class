module example1;
int a;
endmodule
